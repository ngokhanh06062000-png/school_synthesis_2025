//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux_2_1
(
  input  [3:0] d0, d1,
  input        sel,
  output [3:0] y
);

  assign y = sel ? d1 : d0;

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module mux_4_1
(
  input  [3:0] d0, d1, d2, d3,
  input  [1:0] sel,
  output [3:0] y
);

  logic [3:0] low, high;
  mux_2_1 mux_4_1_low(d0, d1, sel[0], low);
  mux_2_1 mux_4_1_high(d2, d3, sel[0], high);
  mux_2_1 mux_4_1_final(low, high, sel[1], y);

endmodule
